.title KiCad schematic
.include "models/BZX84C5V1.spice.txt"
.include "models/C2012C0G2A102J060AA_p.mod"
.include "models/CGJ4C2C0G2A101J060AA_p.mod"
.include "models/FMMT597.spice.txt"
.include "models/SMAZ15.spice.txt"
.include "models/ZXCT1009.spice.txt"
XU4 /SN /PWR_IN /COCM ZXCT1009F
XU5 /PWR_IN /SN CGJ4C2C0G2A101J060AA_p
R6 /SN /PWR_OUT 100
R7 /PWR_IN /PWR_OUT 0.04
R8 /PWR_IN /PWR_OUT 0.04
R5 /SN 0 604k
XU3 /BASE /PWR_IN SMAZ15
R3 0 /BASE 1.5Meg
Q1 /CNV /BASE /COCM FMMT597
R4 /CNV 0 4.99k
R2 /CNV 0 4.99k
R1 /CNV /OUT 100
XU2 /OUT 0 C2012C0G2A102J060AA_p
XU1 0 /OUT DI_BZX84C5V1
V1 /PWR_IN 0 {Vsource}
I1 /PWR_OUT 0 PULSE(0 {Iload} {tdelay} {tr} {tf} {duty} {cycle})
.end
